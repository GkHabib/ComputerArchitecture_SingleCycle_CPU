module TB();

endmodule
