module controller(clk, rst, start, push, pop, memWriteEn, regWriteEn, immAndmem, stm, ldm, branch, jmp, ret, Cin, Zin, opcodeFunc,
  aluOp, cWriteEn, zWriteEn, halt);
